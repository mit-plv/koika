import Complex::*;
import Real::*;
import Vector::*;

import FixedPoint::*;

typedef Complex#(FixedPoint#(16, 16)) ComplexSample;

function ComplexSample getTwiddle(Integer stage, Integer index, Integer points);
    Integer i = ((2*index)/(2 ** (log2(points)-stage))) * (2 ** (log2(points)-stage));
    return cmplx(fromReal(cos(fromInteger(i)*pi/fromInteger(points))),
                 fromReal(-1*sin(fromInteger(i)*pi/fromInteger(points))));
endfunction


module mkGenerate(Empty);
    rule printAll;
        $display("(* Autogenerated by Bluespec\n *)\n");
        $display("Require Import Koika.Frontend.");
        $display("Definition twiddle (stage:nat) (idx:nat) : uaction reg_t ext_fn_t  := match stage, idx with");
   	for(Integer s=0; s<4; s=s+1) begin
		for (Integer i=0; i < 16 ; i=i+1) begin
		let twid = getTwiddle(s,i,16);
		$display("| %d, %d => {{let r := #(Bits.of_N 32 %d) in let i := #(Bits.of_N 32 %d) in struct complex {re:=r;im:=i} }}",s,i, twid.rel,twid.img);
		end
	end
        $display("| _, _ => {{let r := #(Bits.of_N 32 0) in let i := #(Bits.of_N 32 0) in struct complex {re:=r;im:=i} }}");
	$display("end.\n");
	$finish;
    endrule
endmodule

