// -*- verilog -*-
module top(input CLK, input RST_N);
   rv32 core(.CLK, .RST_N);
endmodule

// Local Variables:
// flycheck-verilator-include-path: ("../../_objects/rv32.v/")
// End:
